library ieee;
use ieee.std_logic_1164;
use ieee.numeric_std;

entity robot is 

        generic (

                   n  : integer := 8
        );


end entity;    

